module alu32_tb();
  reg [31:0] A, B;
  reg [2:0] S;
  wire [31:0] R;

  alu32 alu32(A, B, S, R);

  initial begin
    $monitor("%b : %b %b => %b", S, A, B, R);
  end

  initial begin
    #1
      S <= 3'b000; // Add signed
      A <= 128;
      B <= 2;
    #1
      S <= 3'b001; // Sub signed
      A <= 128;
      B <= 2;
    #1
      S <= 3'b010; // And
      A <= 127;
      B <= 2;
    #1
      S <= 3'b011; // Or
      A <= 128;
      B <= 2;
    #1
      S <= 3'b100; // Xor
      A <= 32'b0000_0000_0000_0000_0000_0000_0000_0110;
      B <= 32'b0000_0000_0000_0000_0000_0000_0000_1010;
    #1
      S <= 3'b101; // Sift right arith.
      A <= 32'b1000_0000_0000_0000_0000_0000_0000_1111;
      B <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
    #1
      S <= 3'b110; // Sift right logic
      A <= 32'b1000_0000_0000_0000_0000_0000_0000_1111;
      B <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
    #1
      S <= 3'b111; // Sift left logic
      A <= 32'b1000_0000_0000_0000_0000_0000_0000_1111;
      B <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
  end

endmodule