`include "instDecoder.v"

module instDecoder_tb();

endmodule