`include "module/decoder.v"

module test_decoder();

endmodule