// `include "module/ALU.v"

module ALU_test();
  reg [3:0] i_ctrl;
  reg [31:0] i_1, i_2;
  wire [31:0] o_1;
  wire o_zero, o_neg, o_negU;

  reg [31:0] ans;
  reg res;

  // string op;

  ALU alu(
    .i_ctrl,
    .i_1, .i_2,
    .o_1,
    .o_zero, .o_neg, .o_negU
  );

  // case (i_ctrl)
  //   4'b0000: op = "Add"; 
  //   4': op = ""; 
  //   4': op = ""; 
  //   4': op = ""; 
  //   4': op = ""; 
  //   4': op = ""; 
  //   4': op = ""; 
  //   4': op = ""; 
  //   4': op = ""; 
  //   4': op = ""; 
  //   4': op = ""; 
  //   default: 

  task assert_task;
    #1
    if (o_1 !== ans) begin
      $display("!!!!!!!!!!!!!!!!!!!!!!!!");
      $display("%b failed.", i_ctrl);
      $display("!!!!!!!!!!!!!!!!!!!!!!!!");
      $finish;
    end
  endtask

  // initial begin
  //   $display("++++++++++++++++++++++++");
  //   $display("++++++++++++++++++++++++");
  //   $monitor ("%b(%2d) : %b %b\n", i_ctrl, i_ctrl, i_1, i_2,
  //             "        => %b [z:%b][ng:%b][nU:%b]\n", o_1, o_zero, o_neg, o_negU,
  //             "     ans : %b\n", ans,
  //             "-----------------------");
  // end

  initial begin
        i_1 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        i_2 = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        ans = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
      
    #1
      i_ctrl = 4'b0000; // Add signed
        i_1 = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
        i_2 = 32'b1111_1111_1111_1111_1111_1111_1111_1111;
        ans = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        // assert (o_1 === ans) else $error("0000 Add failed.");
        assert_task;

    #1
      i_ctrl = 4'b0001; // Sub signed
        i_1 = 32'b0000_0000_0000_0000_0000_0000_0000_0100;
        i_2 = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
        ans = 32'b0000_0000_0000_0000_0000_0000_0000_0011;
        assert_task;

    #1
      i_ctrl = 4'b0010; // Or
        i_1 = 32'b0000_0000_0000_0000_0000_0000_0000_0101;
        i_2 = 32'b0000_0000_0000_0000_0000_0000_0000_0011;
        ans = 32'b0000_0000_0000_0000_0000_0000_0000_0111;
        assert_task;

    #1
      i_ctrl = 4'b0011; // And
        i_1 = 32'b0000_0000_0000_0000_0000_0000_0000_0101;
        i_2 = 32'b0000_0000_0000_0000_0000_0000_0000_0011;
        ans = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
        assert_task;

    #1
      i_ctrl = 4'b0100; // Xor
        i_1 = 32'b0000_0000_0000_0000_0000_0000_0000_0101;
        i_2 = 32'b0000_0000_0000_0000_0000_0000_0000_0011;
        ans = 32'b0000_0000_0000_0000_0000_0000_0000_0110;
        assert_task;

    #1
      i_ctrl = 4'b0101; // Sift right arith.
        i_1 = 32'b1000_0000_0000_0000_0000_0000_0000_1111;
        i_2 = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
        ans = 32'b1110_0000_0000_0000_0000_0000_0000_0011;
        assert_task;

    #1
      i_ctrl = 4'b0110; // Sift right logic
        i_1 = 32'b1000_0000_0000_0000_0000_0000_0000_1111;
        i_2 = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
        ans = 32'b0010_0000_0000_0000_0000_0000_0000_0011;
        assert_task;

    #1
      i_ctrl = 4'b0111; // Sift left logic
        i_1 = 32'b1000_0000_0000_0000_0000_0000_0000_1111;
        i_2 = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
        ans = 32'b0000_0000_0000_0000_0000_0000_0011_1100;
        assert_task;

    #1
      i_ctrl = 4'b1101; // Slt
        i_1 = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
        i_2 = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
        ans = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
        assert_task;

      #1
        i_1 = 32'b0000_0000_0000_0000_0000_0000_0000_0100;
        i_2 = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
        ans = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
      #1
        assert_task;

        i_1 = 32'b1000_0000_0000_0000_0000_0000_0000_0000;
        i_2 = 32'b1100_0000_0000_0000_0000_0000_0000_0000;
        ans = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
      #1
        i_1 = 32'b1000_0000_0000_0000_0000_0000_0000_0000;
        i_2 = 32'b0100_0000_0000_0000_0000_0000_0000_0000;
        ans = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
        assert_task;

    #1
      i_ctrl = 4'b1110; // Sltu
        i_1 = 32'b1000_0000_0000_0000_0000_0000_0000_0000;
        i_2 = 32'b0100_0000_0000_0000_0000_0000_0000_0000;
        ans = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        assert_task;

    #1
    $display("assert passed.");
    $finish;
  end
endmodule