module setCause (
  input [3:0] i_causeNum,

  output [3:0] o_cause
);
  assign o_cause = i_causeNum;
  
endmodule